uart/source/uart.vhd